`ifndef __CONFIG_VH__
`define __CONFIG_VH__

`define     BYTEW 8

`define     XADDRW      32
`define     XDATAW      32
`define     XBYTEC      `XDATAW / `BYTEW
`define     XSLAVE_CH   4

`endif