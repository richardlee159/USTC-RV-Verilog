module rom (
    input               xbus_cs,
    input               xbus_we,
    input   [3:0]       xbus_be,
    input   [31:0]      xbus_addr,
    input   [31:0]      xbus_wdata,
    output  [31:0]      xbus_rdata
);

wire [0:63] [31:0] mem  = {
    32'h00000093,
    32'h00000113,
    32'h00000193,
    32'h00000213,
    32'h00000293,
    32'h00000313,
    32'h00000393,
    32'h00000413,
    32'h00000493,
    32'h00000513,
    32'h00000593,
    32'h00000613,
    32'h00000693,
    32'h00000713,
    32'h00000793,
    32'h00000813,
    32'h00000893,
    32'h00000913,
    32'h00000993,
    32'h00000a13,
    32'h00000a93,
    32'h00000b13,
    32'h00000b93,
    32'h00000c13,
    32'h00000c93,
    32'h00000d13,
    32'h00000d93,
    32'h00000e13,
    32'h00000e93,
    32'h00000f13,
    32'h00000f93,
    32'h800000b7,
    32'h00008067
};

wire [5:0] addr = xbus_addr[7:2];

assign xbus_rdata = mem[addr];

endmodule