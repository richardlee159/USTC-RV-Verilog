`ifndef __CONFIG_VH__
`define __CONFIG_VH__

`define NSLAVES 4

`endif